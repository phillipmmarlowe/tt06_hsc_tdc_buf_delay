// This is the unpowered netlist.
module tt_um_hsc_tdc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net16;
 wire net17;
 wire net2;
 wire net3;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \tdc_inst.capt_out[0] ;
 wire \tdc_inst.capt_out[10] ;
 wire \tdc_inst.capt_out[11] ;
 wire \tdc_inst.capt_out[12] ;
 wire \tdc_inst.capt_out[13] ;
 wire \tdc_inst.capt_out[14] ;
 wire \tdc_inst.capt_out[15] ;
 wire \tdc_inst.capt_out[16] ;
 wire \tdc_inst.capt_out[17] ;
 wire \tdc_inst.capt_out[18] ;
 wire \tdc_inst.capt_out[19] ;
 wire \tdc_inst.capt_out[1] ;
 wire \tdc_inst.capt_out[20] ;
 wire \tdc_inst.capt_out[21] ;
 wire \tdc_inst.capt_out[22] ;
 wire \tdc_inst.capt_out[23] ;
 wire \tdc_inst.capt_out[24] ;
 wire \tdc_inst.capt_out[25] ;
 wire \tdc_inst.capt_out[26] ;
 wire \tdc_inst.capt_out[27] ;
 wire \tdc_inst.capt_out[28] ;
 wire \tdc_inst.capt_out[29] ;
 wire \tdc_inst.capt_out[2] ;
 wire \tdc_inst.capt_out[30] ;
 wire \tdc_inst.capt_out[31] ;
 wire \tdc_inst.capt_out[32] ;
 wire \tdc_inst.capt_out[33] ;
 wire \tdc_inst.capt_out[34] ;
 wire \tdc_inst.capt_out[35] ;
 wire \tdc_inst.capt_out[36] ;
 wire \tdc_inst.capt_out[37] ;
 wire \tdc_inst.capt_out[38] ;
 wire \tdc_inst.capt_out[39] ;
 wire \tdc_inst.capt_out[3] ;
 wire \tdc_inst.capt_out[40] ;
 wire \tdc_inst.capt_out[41] ;
 wire \tdc_inst.capt_out[42] ;
 wire \tdc_inst.capt_out[43] ;
 wire \tdc_inst.capt_out[44] ;
 wire \tdc_inst.capt_out[45] ;
 wire \tdc_inst.capt_out[46] ;
 wire \tdc_inst.capt_out[47] ;
 wire \tdc_inst.capt_out[48] ;
 wire \tdc_inst.capt_out[49] ;
 wire \tdc_inst.capt_out[4] ;
 wire \tdc_inst.capt_out[50] ;
 wire \tdc_inst.capt_out[51] ;
 wire \tdc_inst.capt_out[52] ;
 wire \tdc_inst.capt_out[53] ;
 wire \tdc_inst.capt_out[54] ;
 wire \tdc_inst.capt_out[55] ;
 wire \tdc_inst.capt_out[56] ;
 wire \tdc_inst.capt_out[57] ;
 wire \tdc_inst.capt_out[58] ;
 wire \tdc_inst.capt_out[59] ;
 wire \tdc_inst.capt_out[5] ;
 wire \tdc_inst.capt_out[60] ;
 wire \tdc_inst.capt_out[61] ;
 wire \tdc_inst.capt_out[62] ;
 wire \tdc_inst.capt_out[63] ;
 wire \tdc_inst.capt_out[6] ;
 wire \tdc_inst.capt_out[7] ;
 wire \tdc_inst.capt_out[8] ;
 wire \tdc_inst.capt_out[9] ;
 wire \tdc_inst.capt_reg_r[1][0] ;
 wire \tdc_inst.capt_reg_r[1][10] ;
 wire \tdc_inst.capt_reg_r[1][11] ;
 wire \tdc_inst.capt_reg_r[1][12] ;
 wire \tdc_inst.capt_reg_r[1][13] ;
 wire \tdc_inst.capt_reg_r[1][14] ;
 wire \tdc_inst.capt_reg_r[1][15] ;
 wire \tdc_inst.capt_reg_r[1][16] ;
 wire \tdc_inst.capt_reg_r[1][17] ;
 wire \tdc_inst.capt_reg_r[1][18] ;
 wire \tdc_inst.capt_reg_r[1][19] ;
 wire \tdc_inst.capt_reg_r[1][1] ;
 wire \tdc_inst.capt_reg_r[1][20] ;
 wire \tdc_inst.capt_reg_r[1][21] ;
 wire \tdc_inst.capt_reg_r[1][22] ;
 wire \tdc_inst.capt_reg_r[1][23] ;
 wire \tdc_inst.capt_reg_r[1][24] ;
 wire \tdc_inst.capt_reg_r[1][25] ;
 wire \tdc_inst.capt_reg_r[1][26] ;
 wire \tdc_inst.capt_reg_r[1][27] ;
 wire \tdc_inst.capt_reg_r[1][28] ;
 wire \tdc_inst.capt_reg_r[1][29] ;
 wire \tdc_inst.capt_reg_r[1][2] ;
 wire \tdc_inst.capt_reg_r[1][30] ;
 wire \tdc_inst.capt_reg_r[1][31] ;
 wire \tdc_inst.capt_reg_r[1][32] ;
 wire \tdc_inst.capt_reg_r[1][33] ;
 wire \tdc_inst.capt_reg_r[1][34] ;
 wire \tdc_inst.capt_reg_r[1][35] ;
 wire \tdc_inst.capt_reg_r[1][36] ;
 wire \tdc_inst.capt_reg_r[1][37] ;
 wire \tdc_inst.capt_reg_r[1][38] ;
 wire \tdc_inst.capt_reg_r[1][39] ;
 wire \tdc_inst.capt_reg_r[1][3] ;
 wire \tdc_inst.capt_reg_r[1][40] ;
 wire \tdc_inst.capt_reg_r[1][41] ;
 wire \tdc_inst.capt_reg_r[1][42] ;
 wire \tdc_inst.capt_reg_r[1][43] ;
 wire \tdc_inst.capt_reg_r[1][44] ;
 wire \tdc_inst.capt_reg_r[1][45] ;
 wire \tdc_inst.capt_reg_r[1][46] ;
 wire \tdc_inst.capt_reg_r[1][47] ;
 wire \tdc_inst.capt_reg_r[1][48] ;
 wire \tdc_inst.capt_reg_r[1][49] ;
 wire \tdc_inst.capt_reg_r[1][4] ;
 wire \tdc_inst.capt_reg_r[1][50] ;
 wire \tdc_inst.capt_reg_r[1][51] ;
 wire \tdc_inst.capt_reg_r[1][52] ;
 wire \tdc_inst.capt_reg_r[1][53] ;
 wire \tdc_inst.capt_reg_r[1][54] ;
 wire \tdc_inst.capt_reg_r[1][55] ;
 wire \tdc_inst.capt_reg_r[1][56] ;
 wire \tdc_inst.capt_reg_r[1][57] ;
 wire \tdc_inst.capt_reg_r[1][58] ;
 wire \tdc_inst.capt_reg_r[1][59] ;
 wire \tdc_inst.capt_reg_r[1][5] ;
 wire \tdc_inst.capt_reg_r[1][60] ;
 wire \tdc_inst.capt_reg_r[1][61] ;
 wire \tdc_inst.capt_reg_r[1][62] ;
 wire \tdc_inst.capt_reg_r[1][63] ;
 wire \tdc_inst.capt_reg_r[1][6] ;
 wire \tdc_inst.capt_reg_r[1][7] ;
 wire \tdc_inst.capt_reg_r[1][8] ;
 wire \tdc_inst.capt_reg_r[1][9] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[0] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[10] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[11] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[12] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[13] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[14] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[15] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[16] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[17] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[18] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[19] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[1] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[20] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[21] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[22] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[23] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[24] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[25] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[26] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[27] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[28] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[29] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[2] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[30] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[31] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[32] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[33] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[34] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[35] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[36] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[37] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[38] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[39] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[3] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[40] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[41] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[42] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[43] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[44] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[45] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[46] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[47] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[48] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[49] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[4] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[50] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[51] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[52] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[53] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[54] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[55] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[56] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[57] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[58] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[59] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[5] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[60] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[61] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[62] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[63] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[64] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[6] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[7] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[8] ;
 wire \tdc_inst.dl_inst.dl_genblk.dl.ffout_w[9] ;
 wire \tdc_inst.pc_inst.val_in ;
 wire \tdc_inst.pc_inst.val_out ;
 wire \tdc_inst.pg.pg_r_out ;
 wire \tdc_inst.pg.val_r_out ;
 wire \tdc_inst.pg_out ;
 wire \tdc_inst.val_out_capt ;
 wire [1:0] clknet_0_ui_in;
 wire [0:0] clknet_1_0__leaf_ui_in;
 wire [0:0] clknet_1_1__leaf_ui_in;
 wire [1:0] clknet_4_0_0_ui_in;
 wire [1:0] clknet_4_10_0_ui_in;
 wire [1:0] clknet_4_11_0_ui_in;
 wire [1:0] clknet_4_12_0_ui_in;
 wire [1:0] clknet_4_13_0_ui_in;
 wire [1:0] clknet_4_14_0_ui_in;
 wire [1:0] clknet_4_15_0_ui_in;
 wire [1:0] clknet_4_1_0_ui_in;
 wire [1:0] clknet_4_2_0_ui_in;
 wire [1:0] clknet_4_3_0_ui_in;
 wire [1:0] clknet_4_4_0_ui_in;
 wire [1:0] clknet_4_5_0_ui_in;
 wire [1:0] clknet_4_6_0_ui_in;
 wire [1:0] clknet_4_7_0_ui_in;
 wire [1:0] clknet_4_8_0_ui_in;
 wire [1:0] clknet_4_9_0_ui_in;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0077_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__mux2_1 _0469_ (.A0(net151),
    .A1(net6),
    .S(net4),
    .X(_0076_));
 sky130_fd_sc_hd__buf_1 _0470_ (.A(_0076_),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[0] ));
 sky130_fd_sc_hd__inv_2 _0471_ (.A(net12),
    .Y(_0077_));
 sky130_fd_sc_hd__clkbuf_4 _0472_ (.A(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0473_ (.A0(net5),
    .A1(net6),
    .S(net3),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_4 _0474_ (.A(net12),
    .X(_0080_));
 sky130_fd_sc_hd__or2_1 _0475_ (.A(_0080_),
    .B(net151),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_4 _0476_ (.A(net2),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_4 _0477_ (.A(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__o211a_1 _0478_ (.A1(_0078_),
    .A2(_0079_),
    .B1(_0081_),
    .C1(_0083_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_2 _0479_ (.A(_0080_),
    .X(_0084_));
 sky130_fd_sc_hd__or2_1 _0480_ (.A(_0084_),
    .B(net34),
    .X(_0085_));
 sky130_fd_sc_hd__o211a_1 _0481_ (.A1(_0078_),
    .A2(net7),
    .B1(_0083_),
    .C1(_0085_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0482_ (.A0(net34),
    .A1(net7),
    .S(net4),
    .X(_0086_));
 sky130_fd_sc_hd__or2_1 _0483_ (.A(_0080_),
    .B(\tdc_inst.val_out_capt ),
    .X(_0087_));
 sky130_fd_sc_hd__o211a_1 _0484_ (.A1(_0078_),
    .A2(_0086_),
    .B1(_0087_),
    .C1(_0083_),
    .X(_0002_));
 sky130_fd_sc_hd__or2_1 _0485_ (.A(_0084_),
    .B(\tdc_inst.capt_reg_r[1][0] ),
    .X(_0088_));
 sky130_fd_sc_hd__o211a_1 _0486_ (.A1(_0078_),
    .A2(net68),
    .B1(_0083_),
    .C1(_0088_),
    .X(_0003_));
 sky130_fd_sc_hd__or2_1 _0487_ (.A(_0084_),
    .B(\tdc_inst.capt_reg_r[1][1] ),
    .X(_0089_));
 sky130_fd_sc_hd__o211a_1 _0488_ (.A1(_0078_),
    .A2(net72),
    .B1(_0083_),
    .C1(_0089_),
    .X(_0004_));
 sky130_fd_sc_hd__clkbuf_2 _0489_ (.A(_0080_),
    .X(_0090_));
 sky130_fd_sc_hd__or2_1 _0490_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][2] ),
    .X(_0091_));
 sky130_fd_sc_hd__o211a_1 _0491_ (.A1(_0078_),
    .A2(net66),
    .B1(_0083_),
    .C1(_0091_),
    .X(_0005_));
 sky130_fd_sc_hd__buf_2 _0492_ (.A(_0082_),
    .X(_0092_));
 sky130_fd_sc_hd__or2_1 _0493_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][3] ),
    .X(_0093_));
 sky130_fd_sc_hd__o211a_1 _0494_ (.A1(_0078_),
    .A2(net54),
    .B1(_0092_),
    .C1(_0093_),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _0495_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][4] ),
    .X(_0094_));
 sky130_fd_sc_hd__o211a_1 _0496_ (.A1(_0078_),
    .A2(net49),
    .B1(_0092_),
    .C1(_0094_),
    .X(_0007_));
 sky130_fd_sc_hd__or2_1 _0497_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][5] ),
    .X(_0095_));
 sky130_fd_sc_hd__o211a_1 _0498_ (.A1(_0078_),
    .A2(net53),
    .B1(_0092_),
    .C1(_0095_),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _0499_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][6] ),
    .X(_0096_));
 sky130_fd_sc_hd__o211a_1 _0500_ (.A1(_0078_),
    .A2(net99),
    .B1(_0092_),
    .C1(_0096_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _0501_ (.A(_0077_),
    .X(_0097_));
 sky130_fd_sc_hd__or2_1 _0502_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][7] ),
    .X(_0098_));
 sky130_fd_sc_hd__o211a_1 _0503_ (.A1(_0097_),
    .A2(net43),
    .B1(_0092_),
    .C1(_0098_),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _0504_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][8] ),
    .X(_0099_));
 sky130_fd_sc_hd__o211a_1 _0505_ (.A1(_0097_),
    .A2(net51),
    .B1(_0092_),
    .C1(_0099_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _0506_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][9] ),
    .X(_0100_));
 sky130_fd_sc_hd__o211a_1 _0507_ (.A1(_0097_),
    .A2(net82),
    .B1(_0092_),
    .C1(_0100_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _0508_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][10] ),
    .X(_0101_));
 sky130_fd_sc_hd__o211a_1 _0509_ (.A1(_0097_),
    .A2(net39),
    .B1(_0092_),
    .C1(_0101_),
    .X(_0013_));
 sky130_fd_sc_hd__or2_1 _0510_ (.A(_0090_),
    .B(\tdc_inst.capt_reg_r[1][11] ),
    .X(_0102_));
 sky130_fd_sc_hd__o211a_1 _0511_ (.A1(_0097_),
    .A2(net57),
    .B1(_0092_),
    .C1(_0102_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_2 _0512_ (.A(net13),
    .X(_0103_));
 sky130_fd_sc_hd__or2_1 _0513_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][12] ),
    .X(_0104_));
 sky130_fd_sc_hd__o211a_1 _0514_ (.A1(_0097_),
    .A2(net45),
    .B1(_0092_),
    .C1(_0104_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_2 _0515_ (.A(_0082_),
    .X(_0105_));
 sky130_fd_sc_hd__or2_1 _0516_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][13] ),
    .X(_0106_));
 sky130_fd_sc_hd__o211a_1 _0517_ (.A1(_0097_),
    .A2(net62),
    .B1(_0105_),
    .C1(_0106_),
    .X(_0016_));
 sky130_fd_sc_hd__or2_1 _0518_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][14] ),
    .X(_0107_));
 sky130_fd_sc_hd__o211a_1 _0519_ (.A1(_0097_),
    .A2(net46),
    .B1(_0105_),
    .C1(_0107_),
    .X(_0017_));
 sky130_fd_sc_hd__or2_1 _0520_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][15] ),
    .X(_0108_));
 sky130_fd_sc_hd__o211a_1 _0521_ (.A1(_0097_),
    .A2(net47),
    .B1(_0105_),
    .C1(_0108_),
    .X(_0018_));
 sky130_fd_sc_hd__or2_1 _0522_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][16] ),
    .X(_0109_));
 sky130_fd_sc_hd__o211a_1 _0523_ (.A1(_0097_),
    .A2(net97),
    .B1(_0105_),
    .C1(_0109_),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _0524_ (.A(_0077_),
    .X(_0110_));
 sky130_fd_sc_hd__or2_1 _0525_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][17] ),
    .X(_0111_));
 sky130_fd_sc_hd__o211a_1 _0526_ (.A1(_0110_),
    .A2(net74),
    .B1(_0105_),
    .C1(_0111_),
    .X(_0020_));
 sky130_fd_sc_hd__or2_1 _0527_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][18] ),
    .X(_0112_));
 sky130_fd_sc_hd__o211a_1 _0528_ (.A1(_0110_),
    .A2(net105),
    .B1(_0105_),
    .C1(_0112_),
    .X(_0021_));
 sky130_fd_sc_hd__or2_1 _0529_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][19] ),
    .X(_0113_));
 sky130_fd_sc_hd__o211a_1 _0530_ (.A1(_0110_),
    .A2(net123),
    .B1(_0105_),
    .C1(_0113_),
    .X(_0022_));
 sky130_fd_sc_hd__or2_1 _0531_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][20] ),
    .X(_0114_));
 sky130_fd_sc_hd__o211a_1 _0532_ (.A1(_0110_),
    .A2(net78),
    .B1(_0105_),
    .C1(_0114_),
    .X(_0023_));
 sky130_fd_sc_hd__or2_1 _0533_ (.A(_0103_),
    .B(\tdc_inst.capt_reg_r[1][21] ),
    .X(_0115_));
 sky130_fd_sc_hd__o211a_1 _0534_ (.A1(_0110_),
    .A2(net89),
    .B1(_0105_),
    .C1(_0115_),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_2 _0535_ (.A(net17),
    .X(_0116_));
 sky130_fd_sc_hd__or2_1 _0536_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][22] ),
    .X(_0117_));
 sky130_fd_sc_hd__o211a_1 _0537_ (.A1(_0110_),
    .A2(net133),
    .B1(_0105_),
    .C1(_0117_),
    .X(_0025_));
 sky130_fd_sc_hd__buf_2 _0538_ (.A(_0082_),
    .X(_0118_));
 sky130_fd_sc_hd__or2_1 _0539_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][23] ),
    .X(_0119_));
 sky130_fd_sc_hd__o211a_1 _0540_ (.A1(_0110_),
    .A2(net135),
    .B1(_0118_),
    .C1(_0119_),
    .X(_0026_));
 sky130_fd_sc_hd__or2_1 _0541_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][24] ),
    .X(_0120_));
 sky130_fd_sc_hd__o211a_1 _0542_ (.A1(_0110_),
    .A2(net129),
    .B1(_0118_),
    .C1(_0120_),
    .X(_0027_));
 sky130_fd_sc_hd__or2_1 _0543_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][25] ),
    .X(_0121_));
 sky130_fd_sc_hd__o211a_1 _0544_ (.A1(_0110_),
    .A2(net91),
    .B1(_0118_),
    .C1(_0121_),
    .X(_0028_));
 sky130_fd_sc_hd__or2_1 _0545_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][26] ),
    .X(_0122_));
 sky130_fd_sc_hd__o211a_1 _0546_ (.A1(_0110_),
    .A2(net143),
    .B1(_0118_),
    .C1(_0122_),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_4 _0547_ (.A(_0077_),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _0548_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][27] ),
    .X(_0124_));
 sky130_fd_sc_hd__o211a_1 _0549_ (.A1(_0123_),
    .A2(net93),
    .B1(_0118_),
    .C1(_0124_),
    .X(_0030_));
 sky130_fd_sc_hd__or2_1 _0550_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][28] ),
    .X(_0125_));
 sky130_fd_sc_hd__o211a_1 _0551_ (.A1(_0123_),
    .A2(net115),
    .B1(_0118_),
    .C1(_0125_),
    .X(_0031_));
 sky130_fd_sc_hd__or2_1 _0552_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][29] ),
    .X(_0126_));
 sky130_fd_sc_hd__o211a_1 _0553_ (.A1(_0123_),
    .A2(net102),
    .B1(_0118_),
    .C1(_0126_),
    .X(_0032_));
 sky130_fd_sc_hd__or2_1 _0554_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][30] ),
    .X(_0127_));
 sky130_fd_sc_hd__o211a_1 _0555_ (.A1(_0123_),
    .A2(net142),
    .B1(_0118_),
    .C1(_0127_),
    .X(_0033_));
 sky130_fd_sc_hd__or2_1 _0556_ (.A(_0116_),
    .B(\tdc_inst.capt_reg_r[1][31] ),
    .X(_0128_));
 sky130_fd_sc_hd__o211a_1 _0557_ (.A1(_0123_),
    .A2(net36),
    .B1(_0118_),
    .C1(_0128_),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_2 _0558_ (.A(net10),
    .X(_0129_));
 sky130_fd_sc_hd__or2_1 _0559_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][32] ),
    .X(_0130_));
 sky130_fd_sc_hd__o211a_1 _0560_ (.A1(_0123_),
    .A2(net80),
    .B1(_0118_),
    .C1(_0130_),
    .X(_0035_));
 sky130_fd_sc_hd__buf_2 _0561_ (.A(net2),
    .X(_0131_));
 sky130_fd_sc_hd__or2_1 _0562_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][33] ),
    .X(_0132_));
 sky130_fd_sc_hd__o211a_1 _0563_ (.A1(_0123_),
    .A2(net109),
    .B1(_0131_),
    .C1(_0132_),
    .X(_0036_));
 sky130_fd_sc_hd__or2_1 _0564_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][34] ),
    .X(_0133_));
 sky130_fd_sc_hd__o211a_1 _0565_ (.A1(_0123_),
    .A2(net76),
    .B1(_0131_),
    .C1(_0133_),
    .X(_0037_));
 sky130_fd_sc_hd__or2_1 _0566_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][35] ),
    .X(_0134_));
 sky130_fd_sc_hd__o211a_1 _0567_ (.A1(_0123_),
    .A2(net56),
    .B1(_0131_),
    .C1(_0134_),
    .X(_0038_));
 sky130_fd_sc_hd__or2_1 _0568_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][36] ),
    .X(_0135_));
 sky130_fd_sc_hd__o211a_1 _0569_ (.A1(_0123_),
    .A2(net101),
    .B1(_0131_),
    .C1(_0135_),
    .X(_0039_));
 sky130_fd_sc_hd__buf_2 _0570_ (.A(_0077_),
    .X(_0136_));
 sky130_fd_sc_hd__or2_1 _0571_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][37] ),
    .X(_0137_));
 sky130_fd_sc_hd__o211a_1 _0572_ (.A1(_0136_),
    .A2(net149),
    .B1(_0131_),
    .C1(_0137_),
    .X(_0040_));
 sky130_fd_sc_hd__or2_1 _0573_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][38] ),
    .X(_0138_));
 sky130_fd_sc_hd__o211a_1 _0574_ (.A1(_0136_),
    .A2(net131),
    .B1(_0131_),
    .C1(_0138_),
    .X(_0041_));
 sky130_fd_sc_hd__or2_1 _0575_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][39] ),
    .X(_0139_));
 sky130_fd_sc_hd__o211a_1 _0576_ (.A1(_0136_),
    .A2(net126),
    .B1(_0131_),
    .C1(_0139_),
    .X(_0042_));
 sky130_fd_sc_hd__or2_1 _0577_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][40] ),
    .X(_0140_));
 sky130_fd_sc_hd__o211a_1 _0578_ (.A1(_0136_),
    .A2(net59),
    .B1(_0131_),
    .C1(_0140_),
    .X(_0043_));
 sky130_fd_sc_hd__or2_1 _0579_ (.A(_0129_),
    .B(\tdc_inst.capt_reg_r[1][41] ),
    .X(_0141_));
 sky130_fd_sc_hd__o211a_1 _0580_ (.A1(_0136_),
    .A2(net64),
    .B1(_0131_),
    .C1(_0141_),
    .X(_0044_));
 sky130_fd_sc_hd__clkbuf_2 _0581_ (.A(net9),
    .X(_0142_));
 sky130_fd_sc_hd__or2_1 _0582_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][42] ),
    .X(_0143_));
 sky130_fd_sc_hd__o211a_1 _0583_ (.A1(_0136_),
    .A2(net70),
    .B1(_0131_),
    .C1(_0143_),
    .X(_0045_));
 sky130_fd_sc_hd__buf_2 _0584_ (.A(net2),
    .X(_0144_));
 sky130_fd_sc_hd__or2_1 _0585_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][43] ),
    .X(_0145_));
 sky130_fd_sc_hd__o211a_1 _0586_ (.A1(_0136_),
    .A2(net41),
    .B1(_0144_),
    .C1(_0145_),
    .X(_0046_));
 sky130_fd_sc_hd__or2_1 _0587_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][44] ),
    .X(_0146_));
 sky130_fd_sc_hd__o211a_1 _0588_ (.A1(_0136_),
    .A2(net38),
    .B1(_0144_),
    .C1(_0146_),
    .X(_0047_));
 sky130_fd_sc_hd__or2_1 _0589_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][45] ),
    .X(_0147_));
 sky130_fd_sc_hd__o211a_1 _0590_ (.A1(_0136_),
    .A2(net125),
    .B1(_0144_),
    .C1(_0147_),
    .X(_0048_));
 sky130_fd_sc_hd__or2_1 _0591_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][46] ),
    .X(_0148_));
 sky130_fd_sc_hd__o211a_1 _0592_ (.A1(_0136_),
    .A2(net85),
    .B1(_0144_),
    .C1(_0148_),
    .X(_0049_));
 sky130_fd_sc_hd__buf_2 _0593_ (.A(_0077_),
    .X(_0149_));
 sky130_fd_sc_hd__or2_1 _0594_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][47] ),
    .X(_0150_));
 sky130_fd_sc_hd__o211a_1 _0595_ (.A1(_0149_),
    .A2(net145),
    .B1(_0144_),
    .C1(_0150_),
    .X(_0050_));
 sky130_fd_sc_hd__or2_1 _0596_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][48] ),
    .X(_0151_));
 sky130_fd_sc_hd__o211a_1 _0597_ (.A1(_0149_),
    .A2(net121),
    .B1(_0144_),
    .C1(_0151_),
    .X(_0051_));
 sky130_fd_sc_hd__or2_1 _0598_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][49] ),
    .X(_0152_));
 sky130_fd_sc_hd__o211a_1 _0599_ (.A1(_0149_),
    .A2(net147),
    .B1(_0144_),
    .C1(_0152_),
    .X(_0052_));
 sky130_fd_sc_hd__or2_1 _0600_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][50] ),
    .X(_0153_));
 sky130_fd_sc_hd__o211a_1 _0601_ (.A1(_0149_),
    .A2(net119),
    .B1(_0144_),
    .C1(_0153_),
    .X(_0053_));
 sky130_fd_sc_hd__or2_1 _0602_ (.A(_0142_),
    .B(\tdc_inst.capt_reg_r[1][51] ),
    .X(_0154_));
 sky130_fd_sc_hd__o211a_1 _0603_ (.A1(_0149_),
    .A2(net137),
    .B1(_0144_),
    .C1(_0154_),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_2 _0604_ (.A(net8),
    .X(_0155_));
 sky130_fd_sc_hd__or2_1 _0605_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][52] ),
    .X(_0156_));
 sky130_fd_sc_hd__o211a_1 _0606_ (.A1(_0149_),
    .A2(net60),
    .B1(_0144_),
    .C1(_0156_),
    .X(_0055_));
 sky130_fd_sc_hd__buf_2 _0607_ (.A(net2),
    .X(_0157_));
 sky130_fd_sc_hd__or2_1 _0608_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][53] ),
    .X(_0158_));
 sky130_fd_sc_hd__o211a_1 _0609_ (.A1(_0149_),
    .A2(net87),
    .B1(_0157_),
    .C1(_0158_),
    .X(_0056_));
 sky130_fd_sc_hd__or2_1 _0610_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][54] ),
    .X(_0159_));
 sky130_fd_sc_hd__o211a_1 _0611_ (.A1(_0149_),
    .A2(net83),
    .B1(_0157_),
    .C1(_0159_),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _0612_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][55] ),
    .X(_0160_));
 sky130_fd_sc_hd__o211a_1 _0613_ (.A1(_0149_),
    .A2(net128),
    .B1(_0157_),
    .C1(_0160_),
    .X(_0058_));
 sky130_fd_sc_hd__or2_1 _0614_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][56] ),
    .X(_0161_));
 sky130_fd_sc_hd__o211a_1 _0615_ (.A1(_0149_),
    .A2(net111),
    .B1(_0157_),
    .C1(_0161_),
    .X(_0059_));
 sky130_fd_sc_hd__clkbuf_4 _0616_ (.A(_0077_),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _0617_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][57] ),
    .X(_0163_));
 sky130_fd_sc_hd__o211a_1 _0618_ (.A1(_0162_),
    .A2(net103),
    .B1(_0157_),
    .C1(_0163_),
    .X(_0060_));
 sky130_fd_sc_hd__or2_1 _0619_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][58] ),
    .X(_0164_));
 sky130_fd_sc_hd__o211a_1 _0620_ (.A1(_0162_),
    .A2(net138),
    .B1(_0157_),
    .C1(_0164_),
    .X(_0061_));
 sky130_fd_sc_hd__or2_1 _0621_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][59] ),
    .X(_0165_));
 sky130_fd_sc_hd__o211a_1 _0622_ (.A1(_0162_),
    .A2(net95),
    .B1(_0157_),
    .C1(_0165_),
    .X(_0062_));
 sky130_fd_sc_hd__or2_1 _0623_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][60] ),
    .X(_0166_));
 sky130_fd_sc_hd__o211a_1 _0624_ (.A1(_0162_),
    .A2(net140),
    .B1(_0157_),
    .C1(_0166_),
    .X(_0063_));
 sky130_fd_sc_hd__or2_1 _0625_ (.A(_0155_),
    .B(\tdc_inst.capt_reg_r[1][61] ),
    .X(_0167_));
 sky130_fd_sc_hd__o211a_1 _0626_ (.A1(_0162_),
    .A2(net113),
    .B1(_0157_),
    .C1(_0167_),
    .X(_0064_));
 sky130_fd_sc_hd__or2_1 _0627_ (.A(_0080_),
    .B(\tdc_inst.capt_reg_r[1][62] ),
    .X(_0168_));
 sky130_fd_sc_hd__o211a_1 _0628_ (.A1(_0162_),
    .A2(net117),
    .B1(_0157_),
    .C1(_0168_),
    .X(_0065_));
 sky130_fd_sc_hd__or2_1 _0629_ (.A(_0080_),
    .B(\tdc_inst.capt_reg_r[1][63] ),
    .X(_0169_));
 sky130_fd_sc_hd__o211a_1 _0630_ (.A1(_0162_),
    .A2(net152),
    .B1(_0082_),
    .C1(_0169_),
    .X(_0066_));
 sky130_fd_sc_hd__or2_1 _0631_ (.A(\tdc_inst.pc_inst.val_in ),
    .B(_0080_),
    .X(_0170_));
 sky130_fd_sc_hd__o211a_1 _0632_ (.A1(_0162_),
    .A2(net107),
    .B1(_0082_),
    .C1(_0170_),
    .X(_0067_));
 sky130_fd_sc_hd__inv_2 _0633_ (.A(\tdc_inst.capt_reg_r[1][60] ),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _0634_ (.A(\tdc_inst.capt_reg_r[1][42] ),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _0635_ (.A(\tdc_inst.capt_reg_r[1][58] ),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _0636_ (.A(\tdc_inst.capt_reg_r[1][53] ),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _0637_ (.A(\tdc_inst.capt_reg_r[1][49] ),
    .Y(_0175_));
 sky130_fd_sc_hd__nand2_1 _0638_ (.A(\tdc_inst.capt_reg_r[1][43] ),
    .B(\tdc_inst.capt_reg_r[1][39] ),
    .Y(_0176_));
 sky130_fd_sc_hd__or2_1 _0639_ (.A(\tdc_inst.capt_reg_r[1][43] ),
    .B(\tdc_inst.capt_reg_r[1][39] ),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _0640_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__xor2_1 _0641_ (.A(\tdc_inst.capt_reg_r[1][63] ),
    .B(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__inv_2 _0642_ (.A(\tdc_inst.capt_reg_r[1][2] ),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_1 _0643_ (.A(\tdc_inst.capt_reg_r[1][22] ),
    .B(\tdc_inst.capt_reg_r[1][18] ),
    .Y(_0181_));
 sky130_fd_sc_hd__or2_1 _0644_ (.A(\tdc_inst.capt_reg_r[1][22] ),
    .B(\tdc_inst.capt_reg_r[1][18] ),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _0645_ (.A(_0181_),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__xor2_1 _0646_ (.A(\tdc_inst.capt_reg_r[1][35] ),
    .B(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__xnor2_1 _0647_ (.A(_0180_),
    .B(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__xor2_1 _0648_ (.A(_0179_),
    .B(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__xor2_1 _0649_ (.A(\tdc_inst.capt_reg_r[1][28] ),
    .B(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__xnor2_1 _0650_ (.A(\tdc_inst.capt_reg_r[1][5] ),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _0651_ (.A(\tdc_inst.capt_reg_r[1][38] ),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _0652_ (.A(\tdc_inst.capt_reg_r[1][26] ),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _0653_ (.A(\tdc_inst.capt_reg_r[1][23] ),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _0654_ (.A(\tdc_inst.capt_reg_r[1][0] ),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _0655_ (.A(\tdc_inst.capt_reg_r[1][6] ),
    .Y(_0193_));
 sky130_fd_sc_hd__xor2_2 _0656_ (.A(\tdc_inst.capt_reg_r[1][8] ),
    .B(\tdc_inst.capt_reg_r[1][4] ),
    .X(_0194_));
 sky130_fd_sc_hd__xnor2_2 _0657_ (.A(\tdc_inst.capt_reg_r[1][14] ),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__xnor2_2 _0658_ (.A(_0193_),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__xnor2_2 _0659_ (.A(_0192_),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__xnor2_1 _0660_ (.A(_0191_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__xnor2_1 _0661_ (.A(_0190_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__xnor2_1 _0662_ (.A(_0189_),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__xor2_1 _0663_ (.A(_0188_),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_1 _0664_ (.A(\tdc_inst.capt_reg_r[1][47] ),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__or2_1 _0665_ (.A(\tdc_inst.capt_reg_r[1][47] ),
    .B(_0201_),
    .X(_0203_));
 sky130_fd_sc_hd__nand2_1 _0666_ (.A(_0202_),
    .B(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__xnor2_1 _0667_ (.A(_0175_),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _0668_ (.A(\tdc_inst.capt_reg_r[1][34] ),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _0669_ (.A(\tdc_inst.capt_reg_r[1][32] ),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_2 _0670_ (.A(\tdc_inst.capt_reg_r[1][7] ),
    .B(\tdc_inst.capt_reg_r[1][3] ),
    .Y(_0208_));
 sky130_fd_sc_hd__or2_1 _0671_ (.A(\tdc_inst.capt_reg_r[1][7] ),
    .B(\tdc_inst.capt_reg_r[1][3] ),
    .X(_0209_));
 sky130_fd_sc_hd__a21o_1 _0672_ (.A1(_0208_),
    .A2(_0209_),
    .B1(\tdc_inst.capt_reg_r[1][1] ),
    .X(_0210_));
 sky130_fd_sc_hd__nand3_2 _0673_ (.A(\tdc_inst.capt_reg_r[1][1] ),
    .B(_0208_),
    .C(_0209_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _0674_ (.A(_0210_),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _0675_ (.A(\tdc_inst.capt_reg_r[1][11] ),
    .Y(_0213_));
 sky130_fd_sc_hd__xor2_2 _0676_ (.A(\tdc_inst.capt_reg_r[1][17] ),
    .B(\tdc_inst.capt_reg_r[1][13] ),
    .X(_0214_));
 sky130_fd_sc_hd__xnor2_2 _0677_ (.A(\tdc_inst.capt_reg_r[1][10] ),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__xnor2_1 _0678_ (.A(_0213_),
    .B(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__or2_1 _0679_ (.A(_0212_),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__nand2_1 _0680_ (.A(_0212_),
    .B(_0216_),
    .Y(_0218_));
 sky130_fd_sc_hd__and2_1 _0681_ (.A(_0217_),
    .B(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(\tdc_inst.capt_reg_r[1][19] ),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(\tdc_inst.capt_reg_r[1][16] ),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(\tdc_inst.capt_reg_r[1][20] ),
    .Y(_0222_));
 sky130_fd_sc_hd__xor2_2 _0685_ (.A(\tdc_inst.capt_reg_r[1][27] ),
    .B(\tdc_inst.capt_reg_r[1][25] ),
    .X(_0223_));
 sky130_fd_sc_hd__xnor2_2 _0686_ (.A(\tdc_inst.capt_reg_r[1][21] ),
    .B(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__xnor2_2 _0687_ (.A(_0222_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__xnor2_2 _0688_ (.A(_0221_),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__xnor2_2 _0689_ (.A(_0220_),
    .B(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__xor2_1 _0690_ (.A(_0219_),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__or2_1 _0691_ (.A(_0207_),
    .B(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_1 _0692_ (.A(_0207_),
    .B(_0228_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _0693_ (.A(_0229_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__xnor2_2 _0694_ (.A(_0206_),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _0695_ (.A(\tdc_inst.capt_reg_r[1][15] ),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _0696_ (.A(\tdc_inst.capt_reg_r[1][33] ),
    .B(\tdc_inst.capt_reg_r[1][31] ),
    .Y(_0234_));
 sky130_fd_sc_hd__or2_1 _0697_ (.A(\tdc_inst.capt_reg_r[1][33] ),
    .B(\tdc_inst.capt_reg_r[1][31] ),
    .X(_0235_));
 sky130_fd_sc_hd__nand2_1 _0698_ (.A(_0234_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__xor2_2 _0699_ (.A(\tdc_inst.capt_reg_r[1][29] ),
    .B(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(\tdc_inst.capt_reg_r[1][24] ),
    .Y(_0238_));
 sky130_fd_sc_hd__xor2_2 _0701_ (.A(\tdc_inst.capt_reg_r[1][44] ),
    .B(\tdc_inst.capt_reg_r[1][40] ),
    .X(_0239_));
 sky130_fd_sc_hd__xnor2_2 _0702_ (.A(\tdc_inst.capt_reg_r[1][36] ),
    .B(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__xnor2_2 _0703_ (.A(_0238_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__xor2_2 _0704_ (.A(_0237_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__xnor2_2 _0705_ (.A(\tdc_inst.capt_reg_r[1][12] ),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__xnor2_2 _0706_ (.A(_0233_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _0707_ (.A(\tdc_inst.capt_reg_r[1][37] ),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _0708_ (.A(\tdc_inst.capt_reg_r[1][41] ),
    .Y(_0246_));
 sky130_fd_sc_hd__xor2_1 _0709_ (.A(\tdc_inst.capt_reg_r[1][50] ),
    .B(\tdc_inst.capt_reg_r[1][48] ),
    .X(_0247_));
 sky130_fd_sc_hd__xnor2_1 _0710_ (.A(\tdc_inst.capt_reg_r[1][46] ),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__xnor2_1 _0711_ (.A(_0246_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__xnor2_1 _0712_ (.A(_0245_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2_1 _0713_ (.A(\tdc_inst.capt_reg_r[1][57] ),
    .B(\tdc_inst.capt_reg_r[1][54] ),
    .Y(_0251_));
 sky130_fd_sc_hd__or2_1 _0714_ (.A(\tdc_inst.capt_reg_r[1][57] ),
    .B(\tdc_inst.capt_reg_r[1][54] ),
    .X(_0252_));
 sky130_fd_sc_hd__nand2_1 _0715_ (.A(_0251_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__xor2_2 _0716_ (.A(\tdc_inst.capt_reg_r[1][52] ),
    .B(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__inv_2 _0717_ (.A(\tdc_inst.capt_reg_r[1][56] ),
    .Y(_0255_));
 sky130_fd_sc_hd__xor2_2 _0718_ (.A(\tdc_inst.capt_reg_r[1][62] ),
    .B(\tdc_inst.capt_reg_r[1][61] ),
    .X(_0256_));
 sky130_fd_sc_hd__xnor2_2 _0719_ (.A(\tdc_inst.capt_reg_r[1][59] ),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__xnor2_2 _0720_ (.A(_0255_),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__xor2_2 _0721_ (.A(_0254_),
    .B(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__xnor2_1 _0722_ (.A(\tdc_inst.capt_reg_r[1][9] ),
    .B(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__xor2_1 _0723_ (.A(_0250_),
    .B(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__xnor2_1 _0724_ (.A(\tdc_inst.capt_reg_r[1][30] ),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__xor2_1 _0725_ (.A(_0244_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__xnor2_1 _0726_ (.A(\tdc_inst.capt_reg_r[1][45] ),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__xor2_1 _0727_ (.A(_0232_),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__xnor2_1 _0728_ (.A(\tdc_inst.capt_reg_r[1][51] ),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__xor2_1 _0729_ (.A(_0205_),
    .B(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__xnor2_1 _0730_ (.A(\tdc_inst.capt_reg_r[1][55] ),
    .B(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__xnor2_1 _0731_ (.A(_0174_),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__xnor2_2 _0732_ (.A(_0173_),
    .B(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__xnor2_2 _0733_ (.A(_0172_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__nor2_1 _0734_ (.A(_0171_),
    .B(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__and2_1 _0735_ (.A(_0171_),
    .B(_0271_),
    .X(_0273_));
 sky130_fd_sc_hd__o21ai_1 _0736_ (.A1(_0272_),
    .A2(_0273_),
    .B1(_0084_),
    .Y(_0274_));
 sky130_fd_sc_hd__o211a_1 _0737_ (.A1(_0084_),
    .A2(uo_out[0]),
    .B1(_0082_),
    .C1(_0274_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _0738_ (.A(\tdc_inst.capt_reg_r[1][28] ),
    .B(_0186_),
    .X(_0275_));
 sky130_fd_sc_hd__a21o_1 _0739_ (.A1(\tdc_inst.capt_reg_r[1][5] ),
    .A2(_0187_),
    .B1(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__o21ai_2 _0740_ (.A1(_0175_),
    .A2(_0204_),
    .B1(_0202_),
    .Y(_0277_));
 sky130_fd_sc_hd__or2_1 _0741_ (.A(_0189_),
    .B(_0199_),
    .X(_0278_));
 sky130_fd_sc_hd__o21a_1 _0742_ (.A1(_0188_),
    .A2(_0200_),
    .B1(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__o21ai_1 _0743_ (.A1(_0206_),
    .A2(_0231_),
    .B1(_0229_),
    .Y(_0280_));
 sky130_fd_sc_hd__a21bo_1 _0744_ (.A1(\tdc_inst.capt_reg_r[1][63] ),
    .A2(_0177_),
    .B1_N(_0176_),
    .X(_0281_));
 sky130_fd_sc_hd__a21bo_1 _0745_ (.A1(\tdc_inst.capt_reg_r[1][35] ),
    .A2(_0182_),
    .B1_N(_0181_),
    .X(_0282_));
 sky130_fd_sc_hd__or2_1 _0746_ (.A(_0180_),
    .B(_0184_),
    .X(_0283_));
 sky130_fd_sc_hd__o21a_1 _0747_ (.A1(_0179_),
    .A2(_0185_),
    .B1(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__xnor2_1 _0748_ (.A(_0282_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__xor2_1 _0749_ (.A(_0281_),
    .B(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__or2_1 _0750_ (.A(_0193_),
    .B(_0195_),
    .X(_0287_));
 sky130_fd_sc_hd__o21ai_2 _0751_ (.A1(_0192_),
    .A2(_0196_),
    .B1(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__o21ai_2 _0752_ (.A1(_0213_),
    .A2(_0215_),
    .B1(_0217_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand2_1 _0753_ (.A(\tdc_inst.capt_reg_r[1][8] ),
    .B(\tdc_inst.capt_reg_r[1][4] ),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_1 _0754_ (.A(\tdc_inst.capt_reg_r[1][14] ),
    .B(_0194_),
    .Y(_0291_));
 sky130_fd_sc_hd__a22oi_4 _0755_ (.A1(_0290_),
    .A2(_0291_),
    .B1(_0208_),
    .B2(_0211_),
    .Y(_0292_));
 sky130_fd_sc_hd__and4_1 _0756_ (.A(_0290_),
    .B(_0291_),
    .C(_0208_),
    .D(_0211_),
    .X(_0293_));
 sky130_fd_sc_hd__nor2_1 _0757_ (.A(_0292_),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__xnor2_2 _0758_ (.A(_0289_),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__xor2_2 _0759_ (.A(_0288_),
    .B(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__or2_1 _0760_ (.A(_0191_),
    .B(_0197_),
    .X(_0297_));
 sky130_fd_sc_hd__o21a_1 _0761_ (.A1(_0190_),
    .A2(_0198_),
    .B1(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__xor2_1 _0762_ (.A(_0296_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__xnor2_1 _0763_ (.A(_0286_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__xnor2_1 _0764_ (.A(_0280_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__xnor2_2 _0765_ (.A(_0279_),
    .B(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__or2_1 _0766_ (.A(_0220_),
    .B(_0226_),
    .X(_0303_));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(_0227_),
    .Y(_0304_));
 sky130_fd_sc_hd__nand2_1 _0768_ (.A(_0219_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__nand2_1 _0769_ (.A(\tdc_inst.capt_reg_r[1][12] ),
    .B(_0242_),
    .Y(_0306_));
 sky130_fd_sc_hd__o21a_1 _0770_ (.A1(_0233_),
    .A2(_0243_),
    .B1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__and2_1 _0771_ (.A(\tdc_inst.capt_reg_r[1][17] ),
    .B(\tdc_inst.capt_reg_r[1][13] ),
    .X(_0308_));
 sky130_fd_sc_hd__a21oi_1 _0772_ (.A1(\tdc_inst.capt_reg_r[1][10] ),
    .A2(_0214_),
    .B1(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__a21boi_1 _0773_ (.A1(\tdc_inst.capt_reg_r[1][29] ),
    .A2(_0235_),
    .B1_N(_0234_),
    .Y(_0310_));
 sky130_fd_sc_hd__and2_1 _0774_ (.A(\tdc_inst.capt_reg_r[1][27] ),
    .B(\tdc_inst.capt_reg_r[1][25] ),
    .X(_0311_));
 sky130_fd_sc_hd__a21oi_1 _0775_ (.A1(\tdc_inst.capt_reg_r[1][21] ),
    .A2(_0223_),
    .B1(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__or2_1 _0776_ (.A(_0310_),
    .B(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _0777_ (.A(_0310_),
    .B(_0312_),
    .Y(_0314_));
 sky130_fd_sc_hd__nand2_1 _0778_ (.A(_0313_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__or2_1 _0779_ (.A(_0222_),
    .B(_0224_),
    .X(_0316_));
 sky130_fd_sc_hd__o21a_1 _0780_ (.A1(_0221_),
    .A2(_0225_),
    .B1(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__xnor2_1 _0781_ (.A(_0315_),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__xnor2_1 _0782_ (.A(_0309_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__xnor2_1 _0783_ (.A(_0307_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__a21o_1 _0784_ (.A1(_0303_),
    .A2(_0305_),
    .B1(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__nand3_1 _0785_ (.A(_0303_),
    .B(_0305_),
    .C(_0320_),
    .Y(_0322_));
 sky130_fd_sc_hd__and2_2 _0786_ (.A(_0321_),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__or2_1 _0787_ (.A(_0238_),
    .B(_0240_),
    .X(_0324_));
 sky130_fd_sc_hd__o21a_1 _0788_ (.A1(_0237_),
    .A2(_0241_),
    .B1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__or2_1 _0789_ (.A(_0246_),
    .B(_0248_),
    .X(_0326_));
 sky130_fd_sc_hd__o21a_1 _0790_ (.A1(_0245_),
    .A2(_0249_),
    .B1(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__and2_1 _0791_ (.A(\tdc_inst.capt_reg_r[1][44] ),
    .B(\tdc_inst.capt_reg_r[1][40] ),
    .X(_0328_));
 sky130_fd_sc_hd__a21oi_2 _0792_ (.A1(\tdc_inst.capt_reg_r[1][36] ),
    .A2(_0239_),
    .B1(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__xor2_2 _0793_ (.A(_0327_),
    .B(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__xnor2_2 _0794_ (.A(_0325_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__a21bo_2 _0795_ (.A1(\tdc_inst.capt_reg_r[1][52] ),
    .A2(_0252_),
    .B1_N(_0251_),
    .X(_0332_));
 sky130_fd_sc_hd__and2_1 _0796_ (.A(\tdc_inst.capt_reg_r[1][50] ),
    .B(\tdc_inst.capt_reg_r[1][48] ),
    .X(_0333_));
 sky130_fd_sc_hd__a21o_2 _0797_ (.A1(\tdc_inst.capt_reg_r[1][46] ),
    .A2(_0247_),
    .B1(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__xor2_4 _0798_ (.A(_0332_),
    .B(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _0799_ (.A(\tdc_inst.capt_reg_r[1][62] ),
    .B(\tdc_inst.capt_reg_r[1][61] ),
    .X(_0336_));
 sky130_fd_sc_hd__a21o_2 _0800_ (.A1(\tdc_inst.capt_reg_r[1][59] ),
    .A2(_0256_),
    .B1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__or2_1 _0801_ (.A(_0255_),
    .B(_0257_),
    .X(_0338_));
 sky130_fd_sc_hd__o21a_2 _0802_ (.A1(_0254_),
    .A2(_0258_),
    .B1(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__xnor2_4 _0803_ (.A(_0337_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__xnor2_2 _0804_ (.A(_0335_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__nand2_1 _0805_ (.A(\tdc_inst.capt_reg_r[1][9] ),
    .B(_0259_),
    .Y(_0342_));
 sky130_fd_sc_hd__o21a_1 _0806_ (.A1(_0250_),
    .A2(_0260_),
    .B1(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__xor2_2 _0807_ (.A(_0341_),
    .B(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__xnor2_2 _0808_ (.A(_0331_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nand2_1 _0809_ (.A(\tdc_inst.capt_reg_r[1][30] ),
    .B(_0261_),
    .Y(_0346_));
 sky130_fd_sc_hd__o21ai_2 _0810_ (.A1(_0244_),
    .A2(_0262_),
    .B1(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__xnor2_2 _0811_ (.A(_0345_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__xnor2_2 _0812_ (.A(_0323_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__nand2_1 _0813_ (.A(\tdc_inst.capt_reg_r[1][45] ),
    .B(_0263_),
    .Y(_0350_));
 sky130_fd_sc_hd__o21ai_2 _0814_ (.A1(_0232_),
    .A2(_0264_),
    .B1(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__xnor2_2 _0815_ (.A(_0349_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__xnor2_2 _0816_ (.A(_0302_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _0817_ (.A(\tdc_inst.capt_reg_r[1][51] ),
    .B(_0265_),
    .Y(_0354_));
 sky130_fd_sc_hd__o21a_1 _0818_ (.A1(_0205_),
    .A2(_0266_),
    .B1(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__xor2_2 _0819_ (.A(_0353_),
    .B(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__xnor2_2 _0820_ (.A(_0277_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__nand2_1 _0821_ (.A(\tdc_inst.capt_reg_r[1][55] ),
    .B(_0267_),
    .Y(_0358_));
 sky130_fd_sc_hd__o21a_1 _0822_ (.A1(_0174_),
    .A2(_0268_),
    .B1(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__xnor2_2 _0823_ (.A(_0357_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__xor2_2 _0824_ (.A(_0276_),
    .B(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__or2_1 _0825_ (.A(_0173_),
    .B(_0269_),
    .X(_0362_));
 sky130_fd_sc_hd__o21a_1 _0826_ (.A1(_0172_),
    .A2(_0270_),
    .B1(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__xor2_1 _0827_ (.A(_0361_),
    .B(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__xor2_1 _0828_ (.A(_0272_),
    .B(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__or2_1 _0829_ (.A(_0080_),
    .B(uo_out[1]),
    .X(_0366_));
 sky130_fd_sc_hd__o211a_1 _0830_ (.A1(_0162_),
    .A2(_0365_),
    .B1(_0366_),
    .C1(_0083_),
    .X(_0069_));
 sky130_fd_sc_hd__or2_1 _0831_ (.A(_0357_),
    .B(_0359_),
    .X(_0367_));
 sky130_fd_sc_hd__or2b_1 _0832_ (.A(_0360_),
    .B_N(_0276_),
    .X(_0368_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(_0284_),
    .Y(_0369_));
 sky130_fd_sc_hd__and2_1 _0834_ (.A(_0281_),
    .B(_0285_),
    .X(_0370_));
 sky130_fd_sc_hd__a21o_1 _0835_ (.A1(_0282_),
    .A2(_0369_),
    .B1(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__or2b_1 _0836_ (.A(_0300_),
    .B_N(_0280_),
    .X(_0372_));
 sky130_fd_sc_hd__or2b_1 _0837_ (.A(_0279_),
    .B_N(_0301_),
    .X(_0373_));
 sky130_fd_sc_hd__nand2_1 _0838_ (.A(_0372_),
    .B(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__nor2_1 _0839_ (.A(_0296_),
    .B(_0298_),
    .Y(_0375_));
 sky130_fd_sc_hd__a21o_1 _0840_ (.A1(_0286_),
    .A2(_0299_),
    .B1(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__o21ai_1 _0841_ (.A1(_0307_),
    .A2(_0319_),
    .B1(_0321_),
    .Y(_0377_));
 sky130_fd_sc_hd__and2b_1 _0842_ (.A_N(_0295_),
    .B(_0288_),
    .X(_0378_));
 sky130_fd_sc_hd__a21oi_1 _0843_ (.A1(_0289_),
    .A2(_0294_),
    .B1(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__xnor2_1 _0844_ (.A(_0292_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__xor2_1 _0845_ (.A(_0377_),
    .B(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__xor2_1 _0846_ (.A(_0376_),
    .B(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__or2_1 _0847_ (.A(_0315_),
    .B(_0317_),
    .X(_0383_));
 sky130_fd_sc_hd__o21ai_1 _0848_ (.A1(_0309_),
    .A2(_0318_),
    .B1(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__and2b_1 _0849_ (.A_N(_0325_),
    .B(_0330_),
    .X(_0385_));
 sky130_fd_sc_hd__o21ba_1 _0850_ (.A1(_0327_),
    .A2(_0329_),
    .B1_N(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__xnor2_1 _0851_ (.A(_0313_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__xnor2_1 _0852_ (.A(_0384_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__nor2_1 _0853_ (.A(_0341_),
    .B(_0343_),
    .Y(_0389_));
 sky130_fd_sc_hd__a21oi_2 _0854_ (.A1(_0331_),
    .A2(_0344_),
    .B1(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__and2_1 _0855_ (.A(_0332_),
    .B(_0334_),
    .X(_0391_));
 sky130_fd_sc_hd__inv_2 _0856_ (.A(_0337_),
    .Y(_0392_));
 sky130_fd_sc_hd__nor2_1 _0857_ (.A(_0392_),
    .B(_0339_),
    .Y(_0393_));
 sky130_fd_sc_hd__nand2_2 _0858_ (.A(_0391_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__or2_1 _0859_ (.A(_0391_),
    .B(_0393_),
    .X(_0395_));
 sky130_fd_sc_hd__a22oi_4 _0860_ (.A1(_0335_),
    .A2(_0340_),
    .B1(_0394_),
    .B2(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__xor2_1 _0861_ (.A(_0390_),
    .B(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__xnor2_1 _0862_ (.A(_0388_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__or2b_1 _0863_ (.A(_0345_),
    .B_N(_0347_),
    .X(_0399_));
 sky130_fd_sc_hd__a21boi_2 _0864_ (.A1(_0323_),
    .A2(_0348_),
    .B1_N(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__xor2_1 _0865_ (.A(_0398_),
    .B(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__xnor2_1 _0866_ (.A(_0382_),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__and2b_1 _0867_ (.A_N(_0349_),
    .B(_0351_),
    .X(_0403_));
 sky130_fd_sc_hd__a21oi_2 _0868_ (.A1(_0302_),
    .A2(_0352_),
    .B1(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__xnor2_1 _0869_ (.A(_0402_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__xor2_1 _0870_ (.A(_0374_),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__nor2_1 _0871_ (.A(_0353_),
    .B(_0355_),
    .Y(_0407_));
 sky130_fd_sc_hd__a21oi_2 _0872_ (.A1(_0277_),
    .A2(_0356_),
    .B1(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__xor2_1 _0873_ (.A(_0406_),
    .B(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__xnor2_1 _0874_ (.A(_0371_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__a21o_1 _0875_ (.A1(_0367_),
    .A2(_0368_),
    .B1(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__nand3_1 _0876_ (.A(_0367_),
    .B(_0368_),
    .C(_0410_),
    .Y(_0412_));
 sky130_fd_sc_hd__and2_1 _0877_ (.A(_0411_),
    .B(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__nor2_1 _0878_ (.A(_0361_),
    .B(_0363_),
    .Y(_0414_));
 sky130_fd_sc_hd__a21o_1 _0879_ (.A1(_0272_),
    .A2(_0364_),
    .B1(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__or2_1 _0880_ (.A(_0413_),
    .B(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__nand2_1 _0881_ (.A(_0413_),
    .B(_0415_),
    .Y(_0417_));
 sky130_fd_sc_hd__and2_1 _0882_ (.A(_0416_),
    .B(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__or2_1 _0883_ (.A(_0080_),
    .B(uo_out[2]),
    .X(_0419_));
 sky130_fd_sc_hd__o211a_1 _0884_ (.A1(_0162_),
    .A2(_0418_),
    .B1(_0419_),
    .C1(_0083_),
    .X(_0070_));
 sky130_fd_sc_hd__or2_1 _0885_ (.A(_0406_),
    .B(_0408_),
    .X(_0420_));
 sky130_fd_sc_hd__nand2_1 _0886_ (.A(_0371_),
    .B(_0409_),
    .Y(_0421_));
 sky130_fd_sc_hd__nand2_1 _0887_ (.A(_0377_),
    .B(_0380_),
    .Y(_0422_));
 sky130_fd_sc_hd__a21bo_1 _0888_ (.A1(_0376_),
    .A2(_0381_),
    .B1_N(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__nand2_1 _0889_ (.A(_0292_),
    .B(_0378_),
    .Y(_0424_));
 sky130_fd_sc_hd__or2b_1 _0890_ (.A(_0387_),
    .B_N(_0384_),
    .X(_0425_));
 sky130_fd_sc_hd__o21a_1 _0891_ (.A1(_0313_),
    .A2(_0386_),
    .B1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__or2_1 _0892_ (.A(_0424_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _0893_ (.A(_0424_),
    .B(_0426_),
    .Y(_0428_));
 sky130_fd_sc_hd__and2_1 _0894_ (.A(_0427_),
    .B(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__nor2_1 _0895_ (.A(_0390_),
    .B(_0396_),
    .Y(_0430_));
 sky130_fd_sc_hd__a21oi_1 _0896_ (.A1(_0388_),
    .A2(_0397_),
    .B1(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__or2_1 _0897_ (.A(_0394_),
    .B(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__nand2_1 _0898_ (.A(_0394_),
    .B(_0431_),
    .Y(_0433_));
 sky130_fd_sc_hd__and2_1 _0899_ (.A(_0432_),
    .B(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__xnor2_1 _0900_ (.A(_0429_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__nor2_1 _0901_ (.A(_0398_),
    .B(_0400_),
    .Y(_0436_));
 sky130_fd_sc_hd__a21oi_1 _0902_ (.A1(_0382_),
    .A2(_0401_),
    .B1(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__xnor2_1 _0903_ (.A(_0435_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__xor2_1 _0904_ (.A(_0423_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__or2b_1 _0905_ (.A(_0405_),
    .B_N(_0374_),
    .X(_0440_));
 sky130_fd_sc_hd__o21a_1 _0906_ (.A1(_0402_),
    .A2(_0404_),
    .B1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__xnor2_1 _0907_ (.A(_0439_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__a21oi_1 _0908_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__and3_1 _0909_ (.A(_0420_),
    .B(_0421_),
    .C(_0442_),
    .X(_0444_));
 sky130_fd_sc_hd__nor2_1 _0910_ (.A(_0443_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__a21oi_1 _0911_ (.A1(_0411_),
    .A2(_0417_),
    .B1(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__a31o_1 _0912_ (.A1(_0411_),
    .A2(_0417_),
    .A3(_0445_),
    .B1(_0077_),
    .X(_0447_));
 sky130_fd_sc_hd__o221a_1 _0913_ (.A1(_0084_),
    .A2(uo_out[3]),
    .B1(_0446_),
    .B2(_0447_),
    .C1(_0083_),
    .X(_0071_));
 sky130_fd_sc_hd__or2_1 _0914_ (.A(_0439_),
    .B(_0441_),
    .X(_0448_));
 sky130_fd_sc_hd__and2b_1 _0915_ (.A_N(_0438_),
    .B(_0423_),
    .X(_0449_));
 sky130_fd_sc_hd__o21bai_1 _0916_ (.A1(_0435_),
    .A2(_0437_),
    .B1_N(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__a21bo_1 _0917_ (.A1(_0429_),
    .A2(_0434_),
    .B1_N(_0432_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(_0432_),
    .A1(_0451_),
    .S(_0427_),
    .X(_0452_));
 sky130_fd_sc_hd__xnor2_1 _0919_ (.A(_0450_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__nor2_1 _0920_ (.A(_0448_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(_0448_),
    .B(_0453_),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_1 _0922_ (.A(_0454_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__a21o_1 _0923_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0442_),
    .X(_0457_));
 sky130_fd_sc_hd__a21oi_1 _0924_ (.A1(_0411_),
    .A2(_0457_),
    .B1(_0444_),
    .Y(_0458_));
 sky130_fd_sc_hd__a31o_1 _0925_ (.A1(_0413_),
    .A2(_0415_),
    .A3(_0445_),
    .B1(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__xnor2_1 _0926_ (.A(_0456_),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__nand2_1 _0927_ (.A(_0084_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__o211a_1 _0928_ (.A1(_0084_),
    .A2(net154),
    .B1(_0082_),
    .C1(_0461_),
    .X(_0072_));
 sky130_fd_sc_hd__and2b_1 _0929_ (.A_N(_0084_),
    .B(uo_out[5]),
    .X(_0462_));
 sky130_fd_sc_hd__o2bb2a_1 _0930_ (.A1_N(_0450_),
    .A2_N(_0452_),
    .B1(_0427_),
    .B2(_0432_),
    .X(_0463_));
 sky130_fd_sc_hd__a21oi_1 _0931_ (.A1(_0456_),
    .A2(_0459_),
    .B1(_0454_),
    .Y(_0464_));
 sky130_fd_sc_hd__o21ai_1 _0932_ (.A1(_0463_),
    .A2(_0464_),
    .B1(_0080_),
    .Y(_0465_));
 sky130_fd_sc_hd__a21oi_1 _0933_ (.A1(_0463_),
    .A2(_0464_),
    .B1(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__o21a_1 _0934_ (.A1(_0462_),
    .A2(_0466_),
    .B1(_0083_),
    .X(_0073_));
 sky130_fd_sc_hd__o211a_1 _0935_ (.A1(_0084_),
    .A2(uo_out[6]),
    .B1(_0082_),
    .C1(_0465_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(\tdc_inst.pc_inst.val_out ),
    .A1(\tdc_inst.pc_inst.val_in ),
    .S(net15),
    .X(_0467_));
 sky130_fd_sc_hd__and2_1 _0937_ (.A(_0082_),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _0938_ (.A(_0468_),
    .X(_0075_));
 sky130_fd_sc_hd__dfxtp_1 _0939_ (.CLK(clknet_1_0__leaf_ui_in[0]),
    .D(_0000_),
    .Q(\tdc_inst.pg.pg_r_out ));
 sky130_fd_sc_hd__dfxtp_1 _0940_ (.CLK(clknet_1_1__leaf_ui_in[0]),
    .D(_0001_),
    .Q(\tdc_inst.pg.val_r_out ));
 sky130_fd_sc_hd__dfxtp_1 _0941_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(net35),
    .Q(\tdc_inst.val_out_capt ));
 sky130_fd_sc_hd__dfxtp_1 _0942_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(net69),
    .Q(\tdc_inst.capt_reg_r[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0943_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net73),
    .Q(\tdc_inst.capt_reg_r[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0944_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net67),
    .Q(\tdc_inst.capt_reg_r[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0945_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net55),
    .Q(\tdc_inst.capt_reg_r[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0946_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net50),
    .Q(\tdc_inst.capt_reg_r[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0947_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0008_),
    .Q(\tdc_inst.capt_reg_r[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0948_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net100),
    .Q(\tdc_inst.capt_reg_r[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0949_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net44),
    .Q(\tdc_inst.capt_reg_r[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0950_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net52),
    .Q(\tdc_inst.capt_reg_r[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0951_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0012_),
    .Q(\tdc_inst.capt_reg_r[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0952_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(net40),
    .Q(\tdc_inst.capt_reg_r[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0953_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(net58),
    .Q(\tdc_inst.capt_reg_r[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0954_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0015_),
    .Q(\tdc_inst.capt_reg_r[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0955_ (.CLK(clknet_4_11_0_ui_in[1]),
    .D(net63),
    .Q(\tdc_inst.capt_reg_r[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0956_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0017_),
    .Q(\tdc_inst.capt_reg_r[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0957_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(net48),
    .Q(\tdc_inst.capt_reg_r[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0958_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net98),
    .Q(\tdc_inst.capt_reg_r[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0959_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net75),
    .Q(\tdc_inst.capt_reg_r[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0960_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net106),
    .Q(\tdc_inst.capt_reg_r[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0961_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(net124),
    .Q(\tdc_inst.capt_reg_r[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0962_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net79),
    .Q(\tdc_inst.capt_reg_r[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0963_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net90),
    .Q(\tdc_inst.capt_reg_r[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0964_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(net134),
    .Q(\tdc_inst.capt_reg_r[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(net136),
    .Q(\tdc_inst.capt_reg_r[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0966_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(net130),
    .Q(\tdc_inst.capt_reg_r[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net92),
    .Q(\tdc_inst.capt_reg_r[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _0968_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(net144),
    .Q(\tdc_inst.capt_reg_r[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _0969_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net94),
    .Q(\tdc_inst.capt_reg_r[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _0970_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(net116),
    .Q(\tdc_inst.capt_reg_r[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _0971_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(_0032_),
    .Q(\tdc_inst.capt_reg_r[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _0972_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0033_),
    .Q(\tdc_inst.capt_reg_r[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _0973_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(net37),
    .Q(\tdc_inst.capt_reg_r[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _0974_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(net81),
    .Q(\tdc_inst.capt_reg_r[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _0975_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(net110),
    .Q(\tdc_inst.capt_reg_r[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _0976_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(net77),
    .Q(\tdc_inst.capt_reg_r[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _0977_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0038_),
    .Q(\tdc_inst.capt_reg_r[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _0978_ (.CLK(clknet_4_3_0_ui_in[1]),
    .D(_0039_),
    .Q(\tdc_inst.capt_reg_r[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _0979_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(net150),
    .Q(\tdc_inst.capt_reg_r[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(net132),
    .Q(\tdc_inst.capt_reg_r[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(net127),
    .Q(\tdc_inst.capt_reg_r[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0043_),
    .Q(\tdc_inst.capt_reg_r[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(net65),
    .Q(\tdc_inst.capt_reg_r[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net71),
    .Q(\tdc_inst.capt_reg_r[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(net42),
    .Q(\tdc_inst.capt_reg_r[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0047_),
    .Q(\tdc_inst.capt_reg_r[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0048_),
    .Q(\tdc_inst.capt_reg_r[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(net86),
    .Q(\tdc_inst.capt_reg_r[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net146),
    .Q(\tdc_inst.capt_reg_r[1][47] ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(net122),
    .Q(\tdc_inst.capt_reg_r[1][48] ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net148),
    .Q(\tdc_inst.capt_reg_r[1][49] ));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net120),
    .Q(\tdc_inst.capt_reg_r[1][50] ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0054_),
    .Q(\tdc_inst.capt_reg_r[1][51] ));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net61),
    .Q(\tdc_inst.capt_reg_r[1][52] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net88),
    .Q(\tdc_inst.capt_reg_r[1][53] ));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net84),
    .Q(\tdc_inst.capt_reg_r[1][54] ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0058_),
    .Q(\tdc_inst.capt_reg_r[1][55] ));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net112),
    .Q(\tdc_inst.capt_reg_r[1][56] ));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net104),
    .Q(\tdc_inst.capt_reg_r[1][57] ));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net139),
    .Q(\tdc_inst.capt_reg_r[1][58] ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net96),
    .Q(\tdc_inst.capt_reg_r[1][59] ));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net141),
    .Q(\tdc_inst.capt_reg_r[1][60] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net114),
    .Q(\tdc_inst.capt_reg_r[1][61] ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net118),
    .Q(\tdc_inst.capt_reg_r[1][62] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(net153),
    .Q(\tdc_inst.capt_reg_r[1][63] ));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(net108),
    .Q(\tdc_inst.pc_inst.val_in ));
 sky130_fd_sc_hd__dfxtp_4 _1007_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0068_),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfxtp_2 _1008_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0069_),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfxtp_4 _1009_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0070_),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfxtp_4 _1010_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0071_),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfxtp_4 _1011_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0072_),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfxtp_2 _1012_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0073_),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_4 _1013_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0074_),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0075_),
    .Q(\tdc_inst.pc_inst.val_out ));
 sky130_fd_sc_hd__buf_2 _1031_ (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[0] ),
    .X(\tdc_inst.pg_out ));
 sky130_fd_sc_hd__clkbuf_4 _1032_ (.A(\tdc_inst.pc_inst.val_out ),
    .X(uo_out[7]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_ui_in[0]  (.A(ui_in[0]),
    .X(clknet_0_ui_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_ui_in[1]  (.A(ui_in[1]),
    .X(clknet_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_ui_in[0]  (.A(clknet_0_ui_in[0]),
    .X(clknet_1_0__leaf_ui_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_ui_in[0]  (.A(clknet_0_ui_in[0]),
    .X(clknet_1_1__leaf_ui_in[0]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_0_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_0_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_10_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_10_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_11_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_11_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_12_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_12_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_13_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_13_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_14_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_14_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_15_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_15_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_1_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_1_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_2_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_2_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_3_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_3_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_4_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_4_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_5_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_5_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_6_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_6_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_7_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_7_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_8_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_8_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_4_9_0_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_9_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net12),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(net12),
    .X(net11));
 sky130_fd_sc_hd__buf_2 fanout12 (.A(net17),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net17),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net17),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net1),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 fanout8 (.A(net12),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 fanout9 (.A(net12),
    .X(net9));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\tdc_inst.pg.val_r_out ),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\tdc_inst.capt_out[7] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\tdc_inst.capt_out[22] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0025_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\tdc_inst.capt_out[23] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0026_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\tdc_inst.capt_out[51] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\tdc_inst.capt_out[58] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0061_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\tdc_inst.capt_out[60] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0063_),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\tdc_inst.capt_out[30] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0010_),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\tdc_inst.capt_out[26] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0029_),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\tdc_inst.capt_out[47] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0050_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\tdc_inst.capt_out[49] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0052_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\tdc_inst.capt_out[37] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0040_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\tdc_inst.pg.pg_r_out ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\tdc_inst.capt_out[63] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\tdc_inst.capt_out[12] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0066_),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(uo_out[4]),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\tdc_inst.capt_out[14] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\tdc_inst.capt_out[15] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0018_),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\tdc_inst.capt_out[4] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0007_),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\tdc_inst.capt_out[8] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0011_),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0002_),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\tdc_inst.capt_out[5] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\tdc_inst.capt_out[3] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0006_),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\tdc_inst.capt_out[35] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\tdc_inst.capt_out[11] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0014_),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\tdc_inst.capt_out[40] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\tdc_inst.capt_out[52] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0055_),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\tdc_inst.capt_out[13] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\tdc_inst.capt_out[31] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0016_),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\tdc_inst.capt_out[41] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0044_),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\tdc_inst.capt_out[2] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0005_),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\tdc_inst.capt_out[0] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0003_),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\tdc_inst.capt_out[42] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0045_),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\tdc_inst.capt_out[1] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0034_),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0004_),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\tdc_inst.capt_out[17] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0020_),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\tdc_inst.capt_out[34] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0037_),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\tdc_inst.capt_out[20] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0023_),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\tdc_inst.capt_out[32] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0035_),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\tdc_inst.capt_out[9] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\tdc_inst.capt_out[44] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\tdc_inst.capt_out[54] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0057_),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\tdc_inst.capt_out[46] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0049_),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\tdc_inst.capt_out[53] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0056_),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\tdc_inst.capt_out[21] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0024_),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\tdc_inst.capt_out[25] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0028_),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\tdc_inst.capt_out[10] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\tdc_inst.capt_out[27] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0030_),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\tdc_inst.capt_out[59] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0062_),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\tdc_inst.capt_out[16] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0019_),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\tdc_inst.capt_out[6] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0009_),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\tdc_inst.capt_out[36] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\tdc_inst.capt_out[29] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0013_),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\tdc_inst.capt_out[57] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0060_),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\tdc_inst.capt_out[18] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0021_),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\tdc_inst.val_out_capt ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0067_),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\tdc_inst.capt_out[33] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0036_),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\tdc_inst.capt_out[56] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0059_),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\tdc_inst.capt_out[43] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\tdc_inst.capt_out[61] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0064_),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\tdc_inst.capt_out[28] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0031_),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\tdc_inst.capt_out[62] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0065_),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\tdc_inst.capt_out[50] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0053_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\tdc_inst.capt_out[48] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0051_),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0046_),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\tdc_inst.capt_out[19] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_0022_),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\tdc_inst.capt_out[45] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\tdc_inst.capt_out[39] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0042_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\tdc_inst.capt_out[55] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\tdc_inst.capt_out[24] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0027_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\tdc_inst.capt_out[38] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0041_),
    .X(net132));
 sky130_fd_sc_hd__buf_1 input1 (.A(ena),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(rst_n),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[0].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[1] ),
    .DE(net16),
    .Q(\tdc_inst.capt_out[0] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[10].DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[11] ),
    .DE(net15),
    .Q(\tdc_inst.capt_out[10] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[11].DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[12] ),
    .DE(net15),
    .Q(\tdc_inst.capt_out[11] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[12].DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[13] ),
    .DE(net15),
    .Q(\tdc_inst.capt_out[12] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[13].DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[14] ),
    .DE(net14),
    .Q(\tdc_inst.capt_out[13] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[14].DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[15] ),
    .DE(net14),
    .Q(\tdc_inst.capt_out[14] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[15].DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[16] ),
    .DE(net14),
    .Q(\tdc_inst.capt_out[15] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[16].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[17] ),
    .DE(net14),
    .Q(\tdc_inst.capt_out[16] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[17].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[18] ),
    .DE(net14),
    .Q(\tdc_inst.capt_out[17] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[18].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[19] ),
    .DE(net14),
    .Q(\tdc_inst.capt_out[18] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[19].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[20] ),
    .DE(net14),
    .Q(\tdc_inst.capt_out[19] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[1].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[2] ),
    .DE(net16),
    .Q(\tdc_inst.capt_out[1] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[20].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[21] ),
    .DE(net14),
    .Q(\tdc_inst.capt_out[20] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[21].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[22] ),
    .DE(net13),
    .Q(\tdc_inst.capt_out[21] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[22].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[23] ),
    .DE(net13),
    .Q(\tdc_inst.capt_out[22] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[23].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[24] ),
    .DE(net13),
    .Q(\tdc_inst.capt_out[23] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[24].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[25] ),
    .DE(net13),
    .Q(\tdc_inst.capt_out[24] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[25].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[26] ),
    .DE(net13),
    .Q(\tdc_inst.capt_out[25] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[26].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[27] ),
    .DE(net13),
    .Q(\tdc_inst.capt_out[26] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[27].DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[28] ),
    .DE(net13),
    .Q(\tdc_inst.capt_out[27] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[28].DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[29] ),
    .DE(net13),
    .Q(\tdc_inst.capt_out[28] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[29].DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[30] ),
    .DE(net13),
    .Q(\tdc_inst.capt_out[29] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[2].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[3] ),
    .DE(net16),
    .Q(\tdc_inst.capt_out[2] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[30].DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[31] ),
    .DE(net10),
    .Q(\tdc_inst.capt_out[30] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[31].DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[32] ),
    .DE(net11),
    .Q(\tdc_inst.capt_out[31] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[32].DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[33] ),
    .DE(net11),
    .Q(\tdc_inst.capt_out[32] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[33].DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[34] ),
    .DE(net11),
    .Q(\tdc_inst.capt_out[33] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[34].DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[35] ),
    .DE(net11),
    .Q(\tdc_inst.capt_out[34] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[35].DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[36] ),
    .DE(net11),
    .Q(\tdc_inst.capt_out[35] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[36].DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[37] ),
    .DE(net11),
    .Q(\tdc_inst.capt_out[36] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[37].DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[38] ),
    .DE(net11),
    .Q(\tdc_inst.capt_out[37] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[38].DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[39] ),
    .DE(net10),
    .Q(\tdc_inst.capt_out[38] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[39].DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[40] ),
    .DE(net10),
    .Q(\tdc_inst.capt_out[39] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[3].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[4] ),
    .DE(net16),
    .Q(\tdc_inst.capt_out[3] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[40].DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[41] ),
    .DE(net10),
    .Q(\tdc_inst.capt_out[40] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[41].DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[42] ),
    .DE(net10),
    .Q(\tdc_inst.capt_out[41] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[42].DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[43] ),
    .DE(net10),
    .Q(\tdc_inst.capt_out[42] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[43].DFE  (.CLK(clknet_4_6_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[44] ),
    .DE(net10),
    .Q(\tdc_inst.capt_out[43] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[44].DFE  (.CLK(clknet_4_6_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[45] ),
    .DE(net10),
    .Q(\tdc_inst.capt_out[44] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[45].DFE  (.CLK(clknet_4_4_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[46] ),
    .DE(net10),
    .Q(\tdc_inst.capt_out[45] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[46].DFE  (.CLK(clknet_4_4_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[47] ),
    .DE(net9),
    .Q(\tdc_inst.capt_out[46] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[47].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[48] ),
    .DE(net9),
    .Q(\tdc_inst.capt_out[47] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[48].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[49] ),
    .DE(net9),
    .Q(\tdc_inst.capt_out[48] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[49].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[50] ),
    .DE(net9),
    .Q(\tdc_inst.capt_out[49] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[4].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[5] ),
    .DE(net15),
    .Q(\tdc_inst.capt_out[4] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[50].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[51] ),
    .DE(net9),
    .Q(\tdc_inst.capt_out[50] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[51].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[52] ),
    .DE(net9),
    .Q(\tdc_inst.capt_out[51] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[52].DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[53] ),
    .DE(net9),
    .Q(\tdc_inst.capt_out[52] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[53].DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[54] ),
    .DE(net9),
    .Q(\tdc_inst.capt_out[53] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[54].DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[55] ),
    .DE(net9),
    .Q(\tdc_inst.capt_out[54] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[55].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[56] ),
    .DE(net8),
    .Q(\tdc_inst.capt_out[55] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[56].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[57] ),
    .DE(net8),
    .Q(\tdc_inst.capt_out[56] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[57].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[58] ),
    .DE(net8),
    .Q(\tdc_inst.capt_out[57] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[58].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[59] ),
    .DE(net8),
    .Q(\tdc_inst.capt_out[58] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[59].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[60] ),
    .DE(net8),
    .Q(\tdc_inst.capt_out[59] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[5].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[6] ),
    .DE(net15),
    .Q(\tdc_inst.capt_out[5] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[60].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[61] ),
    .DE(net8),
    .Q(\tdc_inst.capt_out[60] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[61].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[62] ),
    .DE(net8),
    .Q(\tdc_inst.capt_out[61] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[62].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[63] ),
    .DE(net8),
    .Q(\tdc_inst.capt_out[62] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[63].DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[64] ),
    .DE(net8),
    .Q(\tdc_inst.capt_out[63] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[6].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[7] ),
    .DE(net15),
    .Q(\tdc_inst.capt_out[6] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[7].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[8] ),
    .DE(net15),
    .Q(\tdc_inst.capt_out[7] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[8].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[9] ),
    .DE(net15),
    .Q(\tdc_inst.capt_out[8] ));
 sky130_fd_sc_hd__edfxtp_1 \tdc_inst.dl_capt.capt_genblk[9].DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[10] ),
    .DE(net15),
    .Q(\tdc_inst.capt_out[9] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[0].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[0] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[1] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[10].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[10] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[11] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[11].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[11] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[12] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[12].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[12] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[13] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[13].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[13] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[14] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[14].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[14] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[15] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[15].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[15] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[16] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[16].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[16] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[17] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[17].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[17] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[18] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[18].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[18] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[19] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[19].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[19] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[20] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[1].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[1] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[2] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[20].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[20] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[21] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[21].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[21] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[22] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[22].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[22] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[23] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[23].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[23] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[24] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[24].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[24] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[25] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[25].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[25] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[26] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[26].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[26] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[27] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[27].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[27] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[28] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[28].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[28] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[29] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[29].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[29] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[30] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[2].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[2] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[3] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[30].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[30] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[31] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[31].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[31] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[32] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[32].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[32] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[33] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[33].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[33] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[34] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[34].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[34] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[35] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[35].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[35] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[36] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[36].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[36] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[37] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[37].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[37] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[38] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[38].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[38] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[39] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[39].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[39] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[40] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[3].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[3] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[4] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[40].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[40] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[41] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[41].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[41] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[42] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[42].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[42] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[43] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[43].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[43] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[44] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[44].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[44] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[45] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[45].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[45] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[46] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[46].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[46] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[47] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[47].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[47] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[48] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[48].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[48] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[49] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[49].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[49] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[50] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[4].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[4] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[5] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[50].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[50] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[51] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[51].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[51] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[52] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[52].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[52] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[53] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[53].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[53] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[54] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[54].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[54] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[55] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[55].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[55] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[56] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[56].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[56] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[57] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[57].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[57] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[58] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[58].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[58] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[59] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[59].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[59] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[60] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[5].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[5] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[6] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[60].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[60] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[61] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[61].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[61] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[62] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[62].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[62] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[63] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[63].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[63] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[64] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[6].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[6] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[7] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[7].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[7] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[8] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[8].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[8] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[9] ));
 sky130_fd_sc_hd__buf_1 \tdc_inst.dl_inst.dl_genblk.dl.dbuf_genblk[9].DB  (.A(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[9] ),
    .X(\tdc_inst.dl_inst.dl_genblk.dl.ffout_w[10] ));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_26 (.HI(net26));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_27 (.HI(net27));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_28 (.HI(net28));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_29 (.HI(net29));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_30 (.HI(net30));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_31 (.HI(net31));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_32 (.HI(net32));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_33 (.HI(net33));
 assign uio_oe[0] = net26;
 assign uio_oe[1] = net27;
 assign uio_oe[2] = net28;
 assign uio_oe[3] = net29;
 assign uio_oe[4] = net30;
 assign uio_oe[5] = net31;
 assign uio_oe[6] = net32;
 assign uio_oe[7] = net33;
 assign uio_out[0] = net18;
 assign uio_out[1] = net19;
 assign uio_out[2] = net20;
 assign uio_out[3] = net21;
 assign uio_out[4] = net22;
 assign uio_out[5] = net23;
 assign uio_out[6] = net24;
 assign uio_out[7] = net25;
endmodule

